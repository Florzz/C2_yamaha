** Profile: "SCHEMATIC1-polarizacion"  [ d:\facu\[8610] dise�o de circuitos electr�nicos\yamaha\yamaha-schematic1-polarizacion.sim ] 

** Creating circuit file "yamaha-schematic1-polarizacion.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad_v2\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\yamaha-SCHEMATIC1.net" 


.END
