** Profile: "SCHEMATIC1-se�al"  [ d:\facu\[8610] dise�o de circuitos electr�nicos\yamaha\yamaha-schematic1-se�al.sim ] 

** Creating circuit file "yamaha-schematic1-se�al.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad_v2\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 3m 0 10000 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\yamaha-SCHEMATIC1.net" 


.END
